// Input
`define CFG_IF_WIDTH    128
`define CFG_IF_HEIGHT   128
`define CFG_IF_CHANNEL  3  
`define CFG_IF_BITWIDTH 16 
`define CFG_IF_FRAC_BIT 8  
`define CFG_IF_PORT     27 

// Kernel/weight
`define CFG_K_WIDTH     3  
`define CFG_K_HEIGHT    3  
`define CFG_K_CHANNEL   3  
`define CFG_K_BITWIDTH  8  
`define CFG_K_FRAC_BIT  6  
`define CFG_K_PORT      1  
`define CFG_K_NUM       3  

// Output
`define CFG_OF_WIDTH    128
`define CFG_OF_HEIGHT   128
`define CFG_OF_CHANNEL  3  
`define CFG_OF_BITWIDTH 16 
`define CFG_OF_FRAC_BIT 8  
`define CFG_OF_PORT     1  
`define CFG_OF_NUM      3  